//Conversor Nacifra-Display de 7 segmentos
module Nasete(
		output reg d7, d6, d5, d4, d3, d2, d1,
		input s5, s4, s3, s2, s1
	     );

	//Conversões:
	/*	s’s	    d’s       ~(d's)
		10000	-> 0000110 -> 1111001
		11000	-> 1011011 -> 0100100
		11100	-> 1001111 -> 0110000
		11110	-> 1100110 -> 0011001
		11111	-> 1101101 -> 0010010
		01111	-> 1111101 -> 0000010
		00111	-> 0000111 -> 1111000
		00011	-> 1111111 -> 0000000
		00001	-> 1101111 -> 0010000s
		00000	-> 0111111 -> 1000000
		invalid -> 1111001 -> 0000110
	*/
	
	always @(*)
		//0000 -> 10000 -> 1111001
		if (s5 == 1 & s4 == 0 & s3 == 0 & s2 == 0 & s1 == 0)
		begin
			d7 = 1;
			d6 = 1;
			d5 = 1;
			d4 = 1;
			d3 = 0;
			d2 = 0;
			d1 = 1;
		end
		//0001 -> 11000 -> 0100100
		else if (s5 == 1 & s4 == 1 & s3 == 0 & s2 == 0 & s1 == 0)
		begin
			d7 = 0;
			d6 = 1;
			d5 = 0;
			d4 = 0;
			d3 = 1;
			d2 = 0;
			d1 = 0;
		end
		//0010 -> 11100 -> 0110000
		else if (s5 == 1 & s4 == 1 & s3 == 1 & s2 == 0 & s1 == 0)
		begin
			d7 = 0;
			d6 = 1;
			d5 = 1;
			d4 = 0;
			d3 = 0;
			d2 = 0;
			d1 = 0;
		end
		//0011 -> 11110 -> 0011001
		else if (s5 == 1 & s4 == 1 & s3 == 1 & s2 == 1 & s1 == 0)
		begin
			d7 = 0;
			d6 = 0;
			d5 = 1;
			d4 = 1;
			d3 = 0;
			d2 = 0;
			d1 = 1;
		end
		//0100 -> 11111 -> 0010010
		else if (s5 == 1 & s4 == 1 & s3 == 1 & s2 == 1 & s1 == 1)
		begin
			d7 = 0;
			d6 = 0;
			d5 = 1;
			d4 = 0;
			d3 = 0;
			d2 = 1;
			d1 = 0;
		end
		//0101 -> 01111 -> 0000010
		else if (s5 == 0 & s4 == 1 & s3 == 1 & s2 == 1 & s1 == 1)
		begin
			d7 = 0;
			d6 = 0;
			d5 = 0;
			d4 = 0;
			d3 = 0;
			d2 = 1;
			d1 = 0;
		end
		//0110 -> 00111 -> 1111000
		else if (s5 == 0 & s4 == 0 & s3 == 1 & s2 == 1 & s1 == 1)
		begin
			d7 = 1;
			d6 = 1;
			d5 = 1;
			d4 = 1;
			d3 = 0;
			d2 = 0;
			d1 = 0;
		end
		//0111 -> 00011 -> 0000000
		else if (s5 == 0 & s4 == 0 & s3 == 0 & s2 == 1 & s1 == 1)
		begin
			d7 = 0;
			d6 = 0;
			d5 = 0;
			d4 = 0;
			d3 = 0;
			d2 = 0;
			d1 = 0;
		end
		//1000 ->00001 -> 0010000
		else if (s5 == 0 & s4 == 0 & s3 == 0 & s2 == 0 & s1 == 1)
		begin
			d7 = 0;
			d6 = 0;
			d5 = 1;
			d4 = 0;
			d3 = 0;
			d2 = 0;
			d1 = 0;
		end
		//1001 -> 00000 -> 1000000
		else if (s5 == 0 & s4 == 0 & s3 == 0 & s2 == 0 & s1 == 0)
		begin
			d7 = 1;
			d6 = 0;
			d5 = 0;
			d4 = 0;
			d3 = 0;
			d2 = 0;
			d1 = 0;
		end
		//invalid -> 0000110
		else 
		begin
			d7 = 0;
			d6 = 0;
			d5 = 0;
			d4 = 0;
			d3 = 1;
			d2 = 1;
			d1 = 0;
		end

endmodule
